//
//	This is the main register code
//	The inputs will be mapped to and from this register file
// This inputs include header hash, difficulty, nonce
//

module register_file ();

endmodule

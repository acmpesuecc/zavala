//
// This file contains the permutation module of the SHA-3 implementation
//

module permutation (
	input logic [1599:0] in_pad,
	input logic clk,
	input logic rst,
	input logic [4:0] op_address,
	output logic [1599:0] readout
};

	// theta function
	
	
	// rho function
	
	
	// pi function
	
	
	// chi function
	
	
	// iota function
	
endmodule
